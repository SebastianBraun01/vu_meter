module ROM (
  input i_clk,
  input [7:0] i_addr,
  input i_ren,
  output reg [23:0] o_data
);

  integer i;
  reg [23:0] register [0:255];

  initial begin
    for (i = 0; i < 256; i = i + 1) register[i] = 'b0;

    // Rote Anzeige
    register[0] = 24'b000000000000111100000000;
    register[1] = 24'b000000000000111100000000;
    register[2] = 24'b000000000000111100000000;
    register[3] = 24'b000000000000111100000000;
    register[4] = 24'b000000000000111100000000;
    register[5] = 24'b000000000000111100000000;
    register[6] = 24'b000000000000111100000000;
    register[7] = 24'b000000000000111100000000;
    register[8] = 24'b000000000000111100000000;
    register[9] = 24'b000000000000111100000000;
    register[10] = 24'b000000000000000000000000;
    register[11] = 24'b000000000000000000000000;
    register[12] = 24'b000000000000000000000000;
    register[13] = 24'b000000000000000000000000;
    register[14] = 24'b000000000000000000000000;
    register[15] = 24'b000000000000000000000000;
    register[16] = 24'b000000000000000000000000;
    register[17] = 24'b000000000000000000000000;
    register[18] = 24'b000000000000000000000000;
    register[19] = 24'b000000000000000000000000;

    // Blaue Anzeige
    register[100] = 24'b000000000000000000000000;
    register[101] = 24'b000000000000000000000000;
    register[102] = 24'b000000000000000000000000;
    register[103] = 24'b000000000000000000000000;
    register[104] = 24'b000000000000000000000000;
    register[105] = 24'b000000000000000000000000;
    register[106] = 24'b000000000000000000000000;
    register[107] = 24'b000000000000000000000000;
    register[108] = 24'b000000000000000000000000;
    register[109] = 24'b000000000000000000000000;
    register[110] = 24'b000000000000000000001111;
    register[111] = 24'b000000000000000000001111;
    register[112] = 24'b000000000000000000001111;
    register[113] = 24'b000000000000000000001111;
    register[114] = 24'b000000000000000000001111;
    register[115] = 24'b000000000000000000001111;
    register[116] = 24'b000000000000000000001111;
    register[117] = 24'b000000000000000000001111;
    register[118] = 24'b000000000000000000001111;
    register[119] = 24'b000000000000000000001111;
  end

  always @(posedge i_clk) begin
    if (i_ren == 1) o_data <= register[i_addr];
    else o_data <= 2'bzz;
  end

endmodule
